`define IOB_ROM_SP_HEXFILE "none"
`define IOB_ROM_SP_ADDR_W 10
`define IOB_ROM_SP_DATA_W 32
`define IOB_ROM_SP_MEM_INIT_FILE_INT {HEXFILE, ".hex"}
`define IOB_ROM_SP_VERSION 16'h0081
