`define IOB_R_DATA_W 1
`define IOB_R_RST_VAL {DATA_W{1'b0}}
`define IOB_R_VERSION 16'h0081
