`define IOB_COUNTER_DATA_W 21
`define IOB_COUNTER_RST_VAL {DATA_W{1'b0}}
`define IOB_COUNTER_VERSION 16'h0081
