`define IOB_CLOCK_CLK_PERIOD 10
`define IOB_CLOCK_VERSION 16'h0081
