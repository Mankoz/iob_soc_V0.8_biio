`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_MERGE_ID_W 0
`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_MERGE_LEN_W 0
`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_MERGE_VERSION 16'h0081
