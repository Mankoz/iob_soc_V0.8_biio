`define IOB_REG_E_DATA_W 21
`define IOB_REG_E_RST_VAL {DATA_W{1'b0}}
`define IOB_REG_E_VERSION 16'h0081
