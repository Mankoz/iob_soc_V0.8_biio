`define IOB_CTLS_VERSION 16'h0081
