`define IOB_RAM_T2P_BE_HEXFILE "none"
`define IOB_RAM_T2P_BE_ADDR_W 0
`define IOB_RAM_T2P_BE_DATA_W 0
`define IOB_RAM_T2P_BE_COL_W 8
`define IOB_RAM_T2P_BE_NUM_COL DATA_W / COL_W
`define IOB_RAM_T2P_BE_MEM_NO_READ_ON_WRITE 0
`define IOB_RAM_T2P_BE_VERSION 16'h0081
