`define IOB_PRIO_ENC_W 21
`define IOB_PRIO_ENC_MODE "LOW"
`define IOB_PRIO_ENC_VERSION 16'h0081
