`define IOB_SOC_SIM_AXI_ID_W 4
`define IOB_SOC_SIM_AXI_LEN_W 8
`define IOB_SOC_SIM_AXI_ADDR_W 15
`define IOB_SOC_SIM_AXI_DATA_W 32
`define IOB_SOC_SIM_BAUD 3000000
`define IOB_SOC_SIM_FREQ 100000000
`define IOB_SOC_SIM_SIMULATION 1
`define IOB_SOC_SIM_VERSION 16'h0081
