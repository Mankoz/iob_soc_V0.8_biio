`timescale 1ns / 1ps
`include "iob_soc_syn_conf.vh"

module iob_soc_syn (
);

endmodule
