`define IOB_SYSTEM_TESTER_IOB_VEXRISCV_AXI_ID_W 0
`define IOB_SYSTEM_TESTER_IOB_VEXRISCV_AXI_ADDR_W 0
`define IOB_SYSTEM_TESTER_IOB_VEXRISCV_AXI_DATA_W 0
`define IOB_SYSTEM_TESTER_IOB_VEXRISCV_AXI_LEN_W 0
`define IOB_SYSTEM_TESTER_IOB_VEXRISCV_VERSION 16'h0001
