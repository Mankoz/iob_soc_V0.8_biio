`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_SPLIT_ID_W 0
`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_SPLIT_LEN_W 0
`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_SPLIT_VERSION 16'h0081
