`define IOB_TIMER_CORE_VERSION 16'h0081
