`define IOB_SOC_PBUS_SPLIT_VERSION 16'h0081
