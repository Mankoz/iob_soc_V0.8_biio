`define IOB_UART_CORE_VERSION 16'h0081
