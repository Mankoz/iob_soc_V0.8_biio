`define IOB_XILINX_CLOCK_WIZARD_OUTPUT_PER 0
`define IOB_XILINX_CLOCK_WIZARD_INPUT_PER 0
`define IOB_XILINX_CLOCK_WIZARD_VERSION 16'h0081
