`define IOB_TIMER_CSRS_ADDR_W 4
`define IOB_TIMER_CSRS_DATA_W 32
`define IOB_TIMER_CSRS_WDATA_W 1
`define IOB_TIMER_CSRS_VERSION 16'h0081
