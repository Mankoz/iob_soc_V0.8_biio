`define IOB_IOB2AXIL_AXIL_ADDR_W 21
`define IOB_IOB2AXIL_AXIL_DATA_W 21
`define IOB_IOB2AXIL_ADDR_W 21
`define IOB_IOB2AXIL_DATA_W 21
`define IOB_IOB2AXIL_VERSION 16'h0081
