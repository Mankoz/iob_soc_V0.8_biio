`define IOB_SOC_SYN_VERSION 16'h0081
