`define IOB_SYSTEM_TESTER_ADDR_W 32
`define IOB_SYSTEM_TESTER_DATA_W 32
`define IOB_SYSTEM_TESTER_INIT_MEM 1
`define IOB_SYSTEM_TESTER_MEM_ADDR_W 18
`define IOB_SYSTEM_TESTER_FW_BASEADDR 0
`define IOB_SYSTEM_TESTER_FW_ADDR_W 18
`define IOB_SYSTEM_TESTER_RST_POL 1
`define IOB_SYSTEM_TESTER_BOOTROM_ADDR_W 12
`define IOB_SYSTEM_TESTER_AXI_ID_W 0
`define IOB_SYSTEM_TESTER_AXI_ADDR_W 18
`define IOB_SYSTEM_TESTER_AXI_DATA_W 32
`define IOB_SYSTEM_TESTER_AXI_LEN_W 4
`define IOB_SYSTEM_TESTER_BOOTROM_MEM_HEXFILE "iob_system_tester_bootrom"
`define IOB_SYSTEM_TESTER_EXT_MEM_HEXFILE "iob_system_tester_firmware"
`define IOB_SYSTEM_TESTER_VERSION 16'h0081
