`define IOB_SYSTEM_TESTER_PBUS_SPLIT_VERSION 16'h0081
