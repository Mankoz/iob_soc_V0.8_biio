`define IOB_SYSTEM_TESTER_SYN_VERSION 16'h0081
