`define IOB_UART_CSRS_ADDR_W 3
`define IOB_UART_CSRS_DATA_W 32
`define IOB_UART_CSRS_RST_POL 1
`define IOB_UART_CSRS_VERSION 16'h0081
