`define IOB_FUNCTIONS_VERSION 16'h0081
