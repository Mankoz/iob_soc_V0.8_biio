`define IOB_BOOTROM_DATA_W 32
`define IOB_BOOTROM_ADDR_W 10
`define IOB_BOOTROM_AXI_ID_W 1
`define IOB_BOOTROM_AXI_LEN_W 8
`define IOB_BOOTROM_VERSION 16'h0081
