`define IOB_SOC_IOB_ZYBO_Z7_AXI_ID_W 4
`define IOB_SOC_IOB_ZYBO_Z7_AXI_LEN_W 8
`define IOB_SOC_IOB_ZYBO_Z7_AXI_ADDR_W 20
`define IOB_SOC_IOB_ZYBO_Z7_AXI_DATA_W 32
`define IOB_SOC_IOB_ZYBO_Z7_BAUD 115200
`define IOB_SOC_IOB_ZYBO_Z7_FREQ 100000000
`define IOB_SOC_IOB_ZYBO_Z7_XILINX 1
`define IOB_SOC_IOB_ZYBO_Z7_VERSION 16'h0081
