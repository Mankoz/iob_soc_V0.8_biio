`define IOB_AXI2IOB_ADDR_WIDTH 32
`define IOB_AXI2IOB_DATA_WIDTH 32
`define IOB_AXI2IOB_STRB_WIDTH (DATA_WIDTH / 8)
`define IOB_AXI2IOB_AXI_ID_WIDTH 8
`define IOB_AXI2IOB_VERSION 16'h0081
