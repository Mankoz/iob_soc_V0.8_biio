`timescale 1ns / 1ps
`include "iob_system_tester_syn_conf.vh"

module iob_system_tester_syn (
);

endmodule
