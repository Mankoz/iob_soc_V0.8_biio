`define IOB_REVERSE_DATA_W 21
`define IOB_REVERSE_VERSION 16'h0081
