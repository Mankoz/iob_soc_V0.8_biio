`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_ID_W 0
`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_LEN_W 0
`define IOB_SYSTEM_TESTER_AXI_FULL_XBAR_VERSION 16'h0081
