`define IOB_PRINTF_VERSION 16'h0081
