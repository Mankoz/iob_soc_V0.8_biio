`define IOB_TASKS_VERSION 16'h0081
